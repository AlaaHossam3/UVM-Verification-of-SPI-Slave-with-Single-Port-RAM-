package Wrapper_config_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh";

    class Wrapper_config extends uvm_object;
        `uvm_object_utils(Wrapper_config)

        virtual Wrapper_if wrapper_vif;
        uvm_active_passive_enum wrapper_is_active;

        function new(string name = "Wrapper_config");
            super.new(name);
        endfunction
    endclass
endpackage

package RAM_agent_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
import RAM_seq_item_pkg::*;
import RAM_driver_pkg::*;
import RAM_monitor_pkg::*;
import RAM_sqr_pkg::*;
import RAM_config_pkg::*;

    class RAM_agent extends uvm_agent;
        `uvm_component_utils(RAM_agent)

        RAM_sqr sqr;
        RAM_driver drv;
        RAM_monitor mon;
        RAM_config cfg;
        uvm_analysis_port #(RAM_seq_item) agt_ap;

        function new(string name = "RAM_agent", uvm_component parent = null);
            super.new(name, parent);
        endfunction

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);

            if(!uvm_config_db #(RAM_config)::get(this, "", "RAM_CFG", cfg))
                `uvm_fatal("Build_phase", "Agent-Unable to get configuration object")
            
            if(cfg.ram_is_active == UVM_ACTIVE) begin
                sqr = RAM_sqr::type_id::create("sqr", this);
                drv = RAM_driver::type_id::create("drv", this);
            end

            mon = RAM_monitor::type_id::create("mon", this);
            agt_ap = new("agt_ap", this);
        endfunction

        function void connect_phase(uvm_phase phase);
            super.connect_phase(phase);

            if(cfg.ram_is_active == UVM_ACTIVE) begin
                drv.ram_vif = cfg.ram_vif;
                drv.seq_item_port.connect(sqr.seq_item_export);
            end

            mon.ram_vif = cfg.ram_vif;
            mon.mon_ap.connect(agt_ap);
        endfunction

    endclass
endpackage